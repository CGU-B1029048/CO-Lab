module lab6(
    input [7:0] A, B;
    input Cin;
    input [2:0] S;
    output [7:0] D;
    output Cout;
);

    
    
endmodule